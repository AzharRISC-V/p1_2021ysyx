module v1 ();
    initial begin
        $display("I am v1");
    end

endmodule //v1
