module v4 (clk);
    input clk;

    v5 u_v5(clk);

endmodule //v1