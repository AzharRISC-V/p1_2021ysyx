module v2 ();
    initial begin
        $display("I am v2");
    end

endmodule //v2