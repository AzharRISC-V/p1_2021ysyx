
// ZhengpuShi

// Cache Top Unit
// 为处理64字节不对齐访问而设计的Cache之上的模块。
// 将可能不对齐的访问转换为1~2次cache访问。

`include "defines.v"

module cache_top (
  input   wire                clk,
  input   wire                rst,
  input   wire  [`BUS_64]     i_cache_top_addr,           // 地址
  input   wire  [`BUS_64]     i_cache_top_wdata,          // 写入的数据
  input   wire  [2 : 0]       i_cache_top_bytes,          // 操作的字节数: 0~7表示1~8字节
	input   wire                i_cache_top_op,             // 操作: 0:read, 1:write
	input   wire                i_cache_top_req,            // 请求
  output  reg   [`BUS_64]     o_cache_top_rdata,          // 读出的数据
	output  reg                 o_cache_top_ack,            // 应答

  // cache_rw 接口
  input   wire  [511:0]       i_cache_rw_axi_rdata,
  input   wire                i_cache_rw_axi_ready,
  output  wire                o_cache_rw_axi_valid,
  output  wire                o_cache_rw_axi_op,
  output  wire  [511:0]       o_cache_rw_axi_wdata,
  output  wire  [63:0]        o_cache_rw_axi_addr,
  output  wire  [1:0]         o_cache_rw_axi_size,
  output  wire  [7:0]         o_cache_rw_axi_blks
);

// =============== cache 从机端 ===============

reg   [63 : 0]                o_cache_addr;        // 存储器地址（字节为单位），64字节对齐，低6位为0。
reg   [63 : 0]                o_cache_wdata;       // 要写入的数据
reg   [2  : 0]                o_cache_bytes;       // 字节数
wire                          o_cache_op;          // 操作类型：0读取，1写入
reg                           o_cache_req;         // 请求
wire  [63 : 0]                i_cache_rdata;       // 已读出的数据
reg                           i_cache_ack;         // 应答

assign o_cache_op = i_cache_top_op;

cache Cache(
  .clk                        (clk                        ),
  .rst                        (rst                        ),
	.i_cache_addr               (o_cache_addr               ),
	.i_cache_wdata              (o_cache_wdata              ),
	.i_cache_bytes              (o_cache_bytes              ),
	.i_cache_op                 (o_cache_op                 ),
	.i_cache_req                (o_cache_req                ),
	.o_cache_rdata              (i_cache_rdata              ),
	.o_cache_ack                (i_cache_ack                ),

  .i_cache_rw_axi_ready       (i_cache_rw_axi_ready       ),
  .i_cache_rw_axi_rdata       (i_cache_rw_axi_rdata       ),
  .o_cache_rw_axi_op          (o_cache_rw_axi_op          ),
  .o_cache_rw_axi_valid       (o_cache_rw_axi_valid       ),
  .o_cache_rw_axi_wdata       (o_cache_rw_axi_wdata       ),
  .o_cache_rw_axi_addr        (o_cache_rw_axi_addr        ),
  .o_cache_rw_axi_size        (o_cache_rw_axi_size        ),
  .o_cache_rw_axi_blks        (o_cache_rw_axi_blks        )
);


// =============== 处理跨行问题 ===============

wire  [59:0]                  i_addr_high;                // 输入地址的高60位
wire  [3:0]                   i_addr_4;                   // 输入地址的低4位 (0~15)
wire  [3:0]                   i_bytes_4;                  // 输入字节数扩展为4位

assign i_addr_high = i_cache_top_addr[63:4];
assign i_addr_4 = i_cache_top_addr[3:0];
assign i_bytes_4 = {1'd0, i_cache_top_bytes};

wire                          en_second;                  // 第二次操作使能
wire  [2 : 0]                 bytes[0:1];                 // 字节数
wire  [63: 0]                 addr[0:1];                  // 地址
wire  [63: 0]                 wdata[0:1];                 // 写数据
reg   [63: 0]                 rdata[0:1];                 // 读数据

assign en_second = i_addr_4 + i_bytes_4 < i_addr_4;
assign bytes[0] = en_second ? {4'd15 - i_addr_4}[2:0] : i_cache_top_bytes;
assign bytes[1] = en_second ? {i_addr_4 + i_bytes_4}[2:0] : 0;
assign addr[0] = i_cache_top_addr;
assign addr[1] = {i_addr_high + 60'd1, 4'd0};
assign wdata[0] = i_cache_top_wdata;
assign wdata[1] = i_cache_top_wdata >> (({3'd0,bytes[0]} + 1) << 3);

wire hs_cache = i_cache_ack & o_cache_req;

assign o_cache_addr = (index == 0) ? addr[0] : addr[1];
assign o_cache_bytes = (index == 0) ? bytes[0] : bytes[1];
assign o_cache_wdata = (index == 0) ? wdata[0] : wdata[1];

reg [1:0]   index;      // 操作的序号：0,1表示两个阶段；其余无效
always @(posedge clk) begin
  if (rst) begin
    index <= 0;
    o_cache_req <= 0;
  end
  else begin
    // 发现用户请求
    if (i_cache_top_req) begin
      // 第一次请求
      if (index == 0) begin
        // 发出请求
        if (!hs_cache) begin
          o_cache_req <= 1;
        end
        // 收到回应
        else begin
          o_cache_req <= 0;
          rdata[0] <= i_cache_rdata;
          // 启动第二次请求，或者结束任务
          if (en_second) begin
            index <= 1;
          end
          else begin
            index <= 3;
            o_cache_top_rdata <= i_cache_rdata;
            o_cache_top_ack <= 1;
          end
        end
      end
      // 第二次请求
      else if (index == 1) begin
        // 发出请求
        if (!hs_cache) begin
          o_cache_req <= 1;
        end
        // 收到回应
        else begin
          rdata[1] <= i_cache_rdata;
          o_cache_top_rdata <= rdata[0] + (i_cache_rdata << ((bytes[0] + 1) << 3));
          o_cache_req <= 0;
          o_cache_top_ack <= 1;
          index <= 3;
        end
      end
    end
    // 结束应答
    else begin
      index <= 0;
      o_cache_top_ack <= 0;
    end
  end
end


endmodule
